.param Vin=24
.param Vout=12
.param Vref=12         ; Reference voltage for closed-loop control
.param fs=100k
.param Pout=10
.param Iout={Pout/Vout}
.param DeltaI=0.083
.param DeltaV=0.12
.param R={Vout/Iout}

; Duty Cycle Calculation
.param D={Vout/Vin}
.param T={1/fs}
.param Ton={D*T}
.param Toff={(1-D)*T}

; Inductor and Capacitor Calculation
.param L={(Vin - Vout)*D/(DeltaI*fs)}
.param C={DeltaI/(8*DeltaV*fs)}

; Gate drive voltage and transition times
.param Vdrive=10
.param trise=10n
.param tfall=10n

; Components
V1 N001 0 {Vin}
L1 N002 Vout {L}
C1 Vout 0 {C}
Rload Vout 0 {R}
D1 0 N002 1N4148
M1 N001 N003 N002 N002 IRFZ44N
Vgate N003 N002 PULSE(0 {Vdrive} {trise} {tfall} {trise} {Ton} {T})

; Error Amplifier (Op-Amp for voltage comparison)
X1 N004 N005 N006 opamp      ; Connect error amplifier here

; PI Controller for duty cycle
X2 N006 N007 PIcontroller      ; Connect PI controller here

; Feedback
Vref N004 0 DC {Vref}         ; Reference voltage for feedback
.model D D
.lib C:\Users\ubai\AppData\Local\LTspice\lib\cmp\standard.dio
.model NMOS NMOS
.model PMOS PMOS
.lib C:\Users\ubai\AppData\Local\LTspice\lib\cmp\standard.mos

* DC-DC Buck Converter with Closed-Loop Control
.include OPAMPmodel.txt    ; Include your op-amp model file
.include PIcontroller.txt  ; Include your PI controller model file
.tran 0 1m 0 1u
.backanno
.end
